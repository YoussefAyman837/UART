interface UART_if;
  logic rx;
  logic tx;
  logic clk;
  logic rst_n;
endinterface //UART_if
  
